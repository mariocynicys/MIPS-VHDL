LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.ALL;
USE IEEE.math_real.ALL;

entity LoadUse is
  port (
    clk   : in std_logic;
    rds
  );
end entity;